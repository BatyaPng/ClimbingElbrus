module log(
    input wire [7:0]num,

    output wire log_num
);

assign log_num = num 