module ms_bit(
    input [7:0]num,

    output wire [3:0]msb
);

assign msb = (num & 8'b10000000) == 8'b10000000 ? 7 :
             (num & 8'b01000000) == 8'b01000000 ? 6 :
             (num & 8'b00100000) == 8'b00100000 ? 5 :
             (num & 8'b00010000) == 8'b00010000 ? 4 :
             (num & 8'b00001000) == 8'b00001000 ? 3 :
             (num & 8'b00000100) == 8'b00000100 ? 2 :
             (num & 8'b00000010) == 8'b00000010 ? 1 :
             (num & 8'b00000001) == 8'b00000001 ? 0 :        
             -1;

endmodule