module normalization (
    input  [48:0] mant_mul,
    output [48:0] mant_norm
);
    

    
endmodule