module muliplier (
    input clk, en,
    input [31:0] op1, op2,

    output [63:0] res,
    output val, overflow
);
    


endmodule   